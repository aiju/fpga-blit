module raminter(
	input wire clk
);

endmodule
